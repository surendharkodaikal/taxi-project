class tx_cfg;
	static string testname;
	static mailbox gen2bfm=new();
	static mailbox mon2cov=new();
	static virtual tx_intf wvif;
endclass
