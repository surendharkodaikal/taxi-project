program tx_tb;
	tx_env env;
	initial begin
		env=new();
		env.run();
	end
endprogram
